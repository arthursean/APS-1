module nota(output wire F, input wire A);
nand(F, A, A);
endmodule